module inst_mem(
	//entrada
	input [31:0] pc,
	
	//saida
	output reg [31:0] rd
);

always @(*)
	begin
	
		/*case(pc)
		8'h00: rd = 32'b000011110011_00000_000_00001_0010011;
		8'h04: rd = 32'b000000001001_00000_000_00010_0010011; 
		8'h08: rd = 32'b0000000_00010_00001_000_00010_0110011;
		8'h0c: rd = 32'b0000000_00010_00001_111_00011_0110011;
		8'h10: rd = 32'b0000000_00010_00001_110_00100_0110011;
		8'h14: rd = 32'b0000000_00100_00011_010_00110_0110011;
		8'h18: rd = 32'b0100000_00110_00100_000_00111_0110011;
		default: rd = 32'b000000000000000000000000000000000;*/
		
		case(pc)
		8'h00: rd = 32'b000011110011_00000_000_00001_0010011;
		8'h04: rd = 32'b000000001001_00000_000_00010_0010011; 
		8'h08: rd = 32'b0000000_00010_00001_000_00010_0110011;
		8'h0c: rd = 32'b0000000_00010_00001_111_00011_0110011;
		8'h10: rd = 32'b0000000_00010_00001_110_00100_0110011;
		8'h14: rd = 32'b0000000_00100_00011_010_00110_0110011;
		8'h18: rd = 32'b0100000_00110_00100_000_00111_0110011;
		default: rd = 32'b000000000000000000000000000000000;
 
		endcase
		
	end

endmodule